// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Davide Rossi <davide.rossi@unibo.it>

module ext_tid_gen
  #(
    parameter EXT_TID_WIDTH = 6
    )
   (
    input   logic                       clk_i,
    input   logic                 rst_ni,

    output  logic                 valid_tid_o,
    output  logic [EXT_TID_WIDTH-1:0]	tid_o,

    input   logic                 incr_i,

    input   logic [EXT_TID_WIDTH-1:0]	tid_i,
    input   logic                       release_tid_i
    );

   localparam NB_OUTSND_TRANS = 2**EXT_TID_WIDTH;

   integer        i;

   logic [127:0]      tid_table;
   logic [6:0]        s_tid;

   always_ff @(posedge clk_i, negedge rst_ni)
     begin
  if(rst_ni == 1'b0)
    begin
       for(i=0; i<NB_OUTSND_TRANS; i++)
         begin
      tid_table[i] <= 1'b0;
         end
       for(i=NB_OUTSND_TRANS; i< 128; i++)
         begin
      tid_table[i] <= 1'b1;
         end
    end
  else
    begin

       if(release_tid_i)
         tid_table[tid_i] <= 1'b0;
       else;

       casex(tid_table)

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0 :
     begin
        if(incr_i)
          begin
       tid_table[0] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01 :
     begin
        if(incr_i)
          begin
       tid_table[1]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011 :
     begin
        if(incr_i)
          begin
       tid_table[2]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111 :
     begin
        if(incr_i)
          begin
       tid_table[3] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111 :
     begin
        if(incr_i)
          begin
       tid_table[4] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111 :
     begin
        if(incr_i)
          begin
       tid_table[5] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111 :
     begin
        if(incr_i)
          begin
       tid_table[6] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[7] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[8] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[9] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[10] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[11] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[12] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[13] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[14] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[15] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[16] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[17] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[18] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[19] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[20] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[21] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[22] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[23] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[24] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[25] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[26] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[27] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[28] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[29] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[30] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[31] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[32] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[33]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[34]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[35] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[36] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[37] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[38] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[39] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[40] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[41] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[42] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[43] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[44] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[45] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[46] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[47] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[48] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[49] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[50] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[51] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[52] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[53] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[54] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[55] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[56] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[57] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[58] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[59] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[60] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[61] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[62] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[63] <= 1'b1;
          end
     end

         //BEGIN
         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[64] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[65]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[66]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[67] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[68] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[69] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[70] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[71] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[72] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[73] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[74] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[75] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[76] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[77] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[78] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[79] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[80] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[81] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[82] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[83] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[84] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[85] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[86] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[87] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[88] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[89] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[90] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[91] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[92] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[93] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[94] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[95] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[96] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[97]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[98]<= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[99] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[100] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[101] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[102] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[103] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[104] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[105] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[106] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[107] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[108] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[109] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[110] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[111] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[112] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[113] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[114] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[115] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[116] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[117] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[118] <= 1'b1;
          end
     end

         128'bxxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[119] <= 1'b1;
          end
     end

         128'bxxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[120] <= 1'b1;
          end
     end

         128'bxxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[121] <= 1'b1;
          end
     end

         128'bxxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[122] <= 1'b1;
          end
     end

         128'bxxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[123] <= 1'b1;
          end
     end

         128'bxxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[124] <= 1'b1;
          end
     end

         128'bxx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[125] <= 1'b1;
          end
     end

         128'bx011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[126] <= 1'b1;
          end
     end

         128'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
     begin
        if(incr_i)
          begin
       tid_table[127] <= 1'b1;
          end
     end

         default:
     begin
     end

       endcase

    end
     end

   always_comb
     begin
  casex(tid_table)

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0 :
      begin
         s_tid            = 0;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01 :
      begin
         s_tid            = 1;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011 :
      begin
         s_tid            = 2;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111 :
      begin
         s_tid            = 3;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111 :
      begin
         s_tid            = 4;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111 :
      begin
         s_tid            = 5;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111 :
      begin
         s_tid            = 6;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111 :
      begin
         s_tid            = 7;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111 :
      begin
         s_tid            = 8;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111 :
      begin
         s_tid            = 9;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111 :
      begin
         s_tid            = 10;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111 :
      begin
         s_tid            = 11;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111 :
      begin
         s_tid            = 12;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111 :
      begin
         s_tid            = 13;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111 :
      begin
         s_tid            = 14;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111 :
      begin
         s_tid            = 15;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111 :
      begin
         s_tid            = 16;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111 :
      begin
         s_tid            = 17;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111 :
      begin
         s_tid            = 18;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111 :
      begin
         s_tid            = 19;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 20;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 21;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxxx_xxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 22;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 23;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 24;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 25;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 26;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 27;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 28;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 29;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 30;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 31;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 32;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 33;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 34;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 35;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 36;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 37;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 38;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 39;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 40;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 41;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 42;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 43;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 44;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 45;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 46;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 47;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 48;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 49;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 50;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 51;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 52;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 53;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 54;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 55;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 56;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 57;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 58;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 59;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 60;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 61;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 62;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 63;
         valid_tid_o      = 1'b1;
      end
//begin
    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 64;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 65;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 66;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 67;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 68;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 69;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 70;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 71;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 72;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 73;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 74;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 75;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 76;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 77;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 78;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 79;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 80;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 81;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 82;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 83;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 84;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 85;
         valid_tid_o      = 1'b1;
      end

    128'bxxxxx_xxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 86;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 87;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 88;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 89;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 90;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 91;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 92;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 93;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 94;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 95;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 96;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 97;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 98;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 99;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 100;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 101;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 102;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 103;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 104;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 105;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 106;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 107;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 108;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 109;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 110;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 111;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 112;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 113;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 114;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 115;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 116;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 117;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 118;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 119;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 120;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_xx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 121;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_x011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 122;
         valid_tid_o      = 1'b1;
      end

    128'bxxxx_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 123;
         valid_tid_o      = 1'b1;
      end

    128'bxxx0_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 124;
         valid_tid_o      = 1'b1;
      end

    128'bxx01_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 125;
         valid_tid_o      = 1'b1;
      end

    128'bx011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 126;
         valid_tid_o      = 1'b1;
      end

    128'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
      begin
         s_tid            = 127;
         valid_tid_o      = 1'b1;
      end
    //end
    default :
      begin
         s_tid            = '0;
         valid_tid_o      = 1'b0;
      end

  endcase

     end

   assign tid_o = s_tid[EXT_TID_WIDTH-1:0];

endmodule

